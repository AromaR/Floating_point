--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   22:52:33 03/27/2015
-- Design Name:   
-- Module Name:   C:/Users/hp/Documents/eda/FPD/tb_div.vhd
-- Project Name:  FPD
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: div
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY tb_div IS
END tb_div;
 
ARCHITECTURE behavior OF tb_div IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT div
    PORT(
         a : IN  std_logic_vector(22 downto 0);
         b : IN  std_logic_vector(22 downto 0);
         c : OUT  std_logic_vector(23 downto 0);
         q : OUT  std_logic_vector(46 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal a : std_logic_vector(22 downto 0) := (others => '0');
   signal b : std_logic_vector(22 downto 0) := (others => '0');

 	--Outputs
   signal c : std_logic_vector(23 downto 0);
   signal q : std_logic_vector(46 downto 0);
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
   --constant <clock>_period : time := 100 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: div PORT MAP (
          a => a,
          b => b,
          c => c,
          q => q
        );

   -- Clock process definitions
--   <clock>_process :process
--   begin
--		<clock> <= '0';
--		wait for <clock>_period/2;
--		<clock> <= '1';
--		wait for <clock>_period/2;
--   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
    a<="11100000000000000000000";
		b<="10000000000000000000000";
		wait for 100 ns;
		a<="11111000000000000000000";
		b<="11000000000000000000000";
		wait for 100 ns;
   end process;

END;
